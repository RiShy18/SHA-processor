/*module expo(Op1, Op2, res);
input [31:0] Op1, Op2;
output [31:0] res;

assign res= Op1**Op2

endmodule
